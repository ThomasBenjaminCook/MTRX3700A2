// LCD_IP.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module LCD_IP (
		input  wire       address,     //   avalon_lcd_slave.address
		input  wire       chipselect,  //                   .chipselect
		input  wire       read,        //                   .read
		input  wire       write,       //                   .write
		input  wire [7:0] writedata,   //                   .writedata
		output wire [7:0] readdata,    //                   .readdata
		output wire       waitrequest, //                   .waitrequest
		input  wire       clk,         //                clk.clk
		inout  wire [7:0] LCD_DATA,    // external_interface.DATA
		output wire       LCD_ON,      //                   .ON
		output wire       LCD_BLON,    //                   .BLON
		output wire       LCD_EN,      //                   .EN
		output wire       LCD_RS,      //                   .RS
		output wire       LCD_RW,      //                   .RW
		input  wire       reset        //              reset.reset
	);

	LCD_IP_character_lcd_0 character_lcd_0 (
		.clk         (clk),         //                clk.clk
		.reset       (reset),       //              reset.reset
		.address     (address),     //   avalon_lcd_slave.address
		.chipselect  (chipselect),  //                   .chipselect
		.read        (read),        //                   .read
		.write       (write),       //                   .write
		.writedata   (writedata),   //                   .writedata
		.readdata    (readdata),    //                   .readdata
		.waitrequest (waitrequest), //                   .waitrequest
		.LCD_DATA    (LCD_DATA),    // external_interface.export
		.LCD_ON      (LCD_ON),      //                   .export
		.LCD_BLON    (LCD_BLON),    //                   .export
		.LCD_EN      (LCD_EN),      //                   .export
		.LCD_RS      (LCD_RS),      //                   .export
		.LCD_RW      (LCD_RW)       //                   .export
	);

endmodule
